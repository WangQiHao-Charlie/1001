`ifndef LSU_OPCODES_VH
`define LSU_OPCODES_VH


parameter LSU_LB = 3'b000;
parameter LSU_LH = 3'b001;
parameter LSU_LW = 3'b010;
parameter LSU_LBU = 3'b011;
parameter LSU_LHU = 3'b100;
parameter LSU_SB = 3'b000;
parameter LSU_SH = 3'b001;
parameter LSU_SW = 3'b010;

`endif
