
module ALU (
    ports
);
    
endmodule